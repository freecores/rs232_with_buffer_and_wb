library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity tb_rx is
end tb_rx;

architecture behaviour of tb_rx is

	--component under test
	component rx_func is
	port(	clk, reset, rx_enable : in std_logic;
			rx : in std_logic;
			
			word_width : in std_logic_vector(3 downto 0);
			baud_period : in std_logic_vector(15 downto 0);
			use_parity_bit, parity_type : in std_logic;
			stop_bits : in std_logic_vector(1 downto 0);
			idle_line_lvl : in std_logic;
			
			start_samples : in std_logic_vector(3 downto 0);	--How many correct samples should give a start bit
			line_samples : in std_logic_vector(3 downto 0);		--How many samples should tip the internal rx value
			
			data 		: out std_logic_vector(7 downto 0);
			data_ready 	: out std_logic;
			parity_error :	out std_logic;
			stop_bit_error : out std_logic);
	end component;

	--tx_func is only used for generating signals
	component tx_func is
	port(	clk, reset : in std_logic;
			data : in std_logic_vector(7 downto 0);
			transmit_data : in std_logic;
			
			word_width : in std_logic_vector(3 downto 0);
			baud_period : in std_logic_vector(15 downto 0);
			use_parity_bit, parity_type : in std_logic;
			stop_bits : in std_logic_vector(1 downto 0);
			idle_line_lvl : in std_logic;

			tx : out std_logic;
			sending : out std_logic);
	end component;
	
	
	signal clk : std_logic := '0';
	signal reset : std_logic := '0';	
	constant clk_period : time := 2 ns;	-- 50MHz
	
	signal transmit_data : std_logic := '0';
	signal word_width : std_logic_vector(3 downto 0) := "1000";
	signal baud_period : std_logic_vector(15 downto 0) := "0000000000100000";
	signal use_parity_bit : std_logic := '1';
	signal parity_type : std_logic := '0';	--0 = even, 1 = odd
	signal stop_bits : std_logic_vector(1 downto 0) := "01";

	signal txrx, sending : std_logic;
	signal idle_line_lvl : std_logic := '1';
	
	signal tx_data : std_logic_vector(7 downto 0) := "00000000";
	signal rx_data : std_logic_vector(7 downto 0);

	--specific for rx_func
	signal rx_enable : std_logic := '1';
	signal start_samples : std_logic_vector(3 downto 0) := "1100";	--How many correct samples should give a start bit
	signal line_samples : std_logic_vector(3 downto 0) := "0100";	--How many samples should tip the internal rx value
	signal data_ready : std_logic;
	signal parity_error : std_logic;
	signal stop_bit_error : std_logic;

	signal stimuli_input	: std_logic_vector(7 downto 0) := "00000000";
	signal expected_output 	: std_logic_vector(7 downto 0) := "00000000";

begin

	--unit under test
	uut0 : rx_func port map (clk, reset, rx_enable, txrx, word_width, baud_period, use_parity_bit, parity_type, stop_bits, idle_line_lvl, start_samples, line_samples, rx_data, data_ready, parity_error, stop_bit_error);

	uut1 : tx_func port map (clk, reset, tx_data, transmit_data, word_width, baud_period, use_parity_bit, parity_type, stop_bits, idle_line_lvl, txrx, sending);
	
	clk_process : process
	begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2; 
	end process;
	
	reset_process : process
	begin
		reset <= '0';
		wait for 12 ns;
		reset <= '1';
		wait for 5 ns;
		reset <= '0';
		wait;
	end process;
	
	new_data_process : process
	begin
		wait until reset = '1';
		wait until reset = '0';
		wait for 5 ns;
		tx_data <= "00000000";
		transmit_data <= '1';
		wait for 2 ns;
		transmit_data <= '0';
		
		
		while stimuli_input /= "11111111" loop
			wait until sending = '0';
			wait for 12 ns;

			tx_data <= tx_data + '1';
			transmit_data <= '1';
			wait for 2 ns;
			transmit_data <= '0';
		end loop;
		
		wait;		
	end process;
	
	data_check : process
	begin
		wait until data_ready = '1';
			assert rx_data = expected_output report "Not expected output" severity warning;
		wait until data_ready = '0';
		expected_output <= expected_output + 1;
		
		if expected_output = "11111111" then
			wait until data_ready = '1';
			assert rx_data = expected_output report "Not expected output" severity warning;
			wait until data_ready = '0';
			wait for 100 ns;
			assert false report "None - end of simulation" severity failure;
		end if;
	end process;

	protocol_error : process
	begin
		wait for 1 ns;
		assert parity_error = '0' report "Stob bit error" severity error;
		assert stop_bit_error = '0' report "Stob bit error" severity error;
	end process;
	
end behaviour;